-- $Id: ram32k_b16.vhd,v 1.2 2008/03/14 15:52:43 dilbert57 Exp $
--===========================================================================--
--                                                                           --
--  ram32k_b16.vhd - 32KByte Block RAM Component for Spartan 3/3E            --
--                                                                           --
--===========================================================================--
--
--  File name      : ram32k_b16.vhd
--
--  Entity name    : ram_32k
--
--  Purpose        : Implements 32K of Synchronous Static RAM 
--                   using 16 x Spartan 3/3E RAMB16_S9 block rams
--                   Used in the Digilent Spartan 3E500 System09 design
--                  
--  Dependencies   : ieee.Std_Logic_1164
--                   ieee.std_logic_arith
--                   unisim.vcomponents
--
--  Uses           : RAMB16_S9
--
--  Author         : John E. Kent
--
--  Email          : dilbert57@opencores.org      
--
--  Web            : http://opencores.org/project,system09
--
--
--  Copyright (C) 2005 - 2010 John Kent
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--===========================================================================--
--                                                                           --
--                              Revision  History                            --
--                                                                           --
--===========================================================================--
--
-- Version Author      Date          Changes
--
-- 0.1     John Kent   2006-04-24    Initial release
-- 0.2     John Kent   2005-06-29    Added CS term to CE decodes. (date ???)
-- 0.3     John Kent   2010-09-14    Renamed "rdata" to "data_out"
--                                   Renamed "wdata" to "data_in"
--                                   Added header description
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.vcomponents.all;

entity ram_32k is
    Port (
       clk      : in  std_logic;
		 rst      : in  std_logic;
		 cs       : in  std_logic;
       addr     : in  std_logic_vector (14 downto 0);
		 rw       : in  std_logic;
       data_in  : in  std_logic_vector (7 downto 0);
       data_out : out std_logic_vector (7 downto 0)
    );
end ram_32k;

architecture rtl of ram_32k is


signal we         : std_logic;
signal dp         : std_logic_vector(15 downto 0);
signal ce         : std_logic_vector(15 downto 0);
signal data_out_0 : std_logic_vector(7 downto 0);
signal data_out_1 : std_logic_vector(7 downto 0);
signal data_out_2 : std_logic_vector(7 downto 0);
signal data_out_3 : std_logic_vector(7 downto 0);
signal data_out_4 : std_logic_vector(7 downto 0);
signal data_out_5 : std_logic_vector(7 downto 0);
signal data_out_6 : std_logic_vector(7 downto 0);
signal data_out_7 : std_logic_vector(7 downto 0);
signal data_out_8 : std_logic_vector(7 downto 0);
signal data_out_9 : std_logic_vector(7 downto 0);
signal data_out_a : std_logic_vector(7 downto 0);
signal data_out_b : std_logic_vector(7 downto 0);
signal data_out_c : std_logic_vector(7 downto 0);
signal data_out_d : std_logic_vector(7 downto 0);
signal data_out_e : std_logic_vector(7 downto 0);
signal data_out_f : std_logic_vector(7 downto 0);

begin

  RAM0 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_0,
	  dop(0) => dp(0),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(0),
	  en   => ce(0),
	  ssr  => rst,
	  we   => we
	);

  RAM1 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_1,
	  dop(0) => dp(1),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(1),
	  en   => ce(1),
	  ssr  => rst,
	  we   => we
	);

  RAM2 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_2,
	  dop(0) => dp(2),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(2),
	  en   => ce(2),
	  ssr  => rst,
	  we   => we
	);

  RAM3 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_3,
	  dop(0) => dp(3),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(3),
	  en   => ce(3),
	  ssr  => rst,
	  we   => we
	);

  RAM4 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_4,
	  dop(0) => dp(4),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(4),
	  en   => ce(4),
	  ssr  => rst,
	  we   => we
	);

  RAM5 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_5,
	  dop(0) => dp(5),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(5),
	  en   => ce(5),
	  ssr  => rst,
	  we   => we
	);

  RAM6 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_6,
	  dop(0) => dp(6),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(6),
	  en   => ce(6),
	  ssr  => rst,
	  we   => we
	);

  RAM7 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_7,
	  dop(0) => dp(7),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(7),
	  en   => ce(7),
	  ssr  => rst,
	  we   => we
	);

  RAM8 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_8,
	  dop(0) => dp(8),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(8),
	  en   => ce(8),
	  ssr  => rst,
	  we   => we
	);

  RAM9 : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_9,
	  dop(0) => dp(9),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(9),
	  en   => ce(9),
	  ssr  => rst,
	  we   => we
	);

  RAMA : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_a,
	  dop(0) => dp(10),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(10),
	  en   => ce(10),
	  ssr  => rst,
	  we   => we
	);

  RAMB : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_b,
	  dop(0) => dp(11),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(11),
	  en   => ce(11),
	  ssr  => rst,
	  we   => we
	);

  RAMC : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_c,
	  dop(0) => dp(12),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(12),
	  en   => ce(12),
	  ssr  => rst,
	  we   => we
	);

  RAMD : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_d,
	  dop(0) => dp(13),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(13),
	  en   => ce(13),
	  ssr  => rst,
	  we   => we
	);

  RAME : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_e,
	  dop(0) => dp(14),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(14),
	  en   => ce(14),
	  ssr  => rst,
	  we   => we
	);

  RAMF : RAMB16_S9
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map (
	  do   => data_out_f,
	  dop(0) => dp(15),
	  addr => addr(10 downto 0),
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp(15),
	  en   => ce(15),
	  ssr  => rst,
	  we   => we
	);

my_ram_32k : process ( cs, rw, addr,
                       data_out_0, data_out_1, data_out_2, data_out_3,
                       data_out_4, data_out_5, data_out_6, data_out_7,
                       data_out_8, data_out_9, data_out_a, data_out_b,
                       data_out_c, data_out_d, data_out_e, data_out_f )
begin
	 we <= not rw;
	 
	 case addr(14 downto 11) is
	 when "0000" =>
	     data_out <= data_out_0;
	 when "0001" =>
	     data_out <= data_out_1;
	 when "0010" =>
	     data_out <= data_out_2;
	 when "0011" =>
	     data_out <= data_out_3;
	 when "0100" =>
	     data_out <= data_out_4;
	 when "0101" =>
	     data_out <= data_out_5;
	 when "0110" =>
	     data_out <= data_out_6;
	 when "0111" =>
	     data_out <= data_out_7;
	 when "1000" =>
	     data_out <= data_out_8;
	 when "1001" =>
	     data_out <= data_out_9;
	 when "1010" =>
	     data_out <= data_out_a;
	 when "1011" =>
	     data_out <= data_out_b;
	 when "1100" =>
	     data_out <= data_out_c;
	 when "1101" =>
	     data_out <= data_out_d;
	 when "1110" =>
	     data_out <= data_out_e;
	 when "1111" =>
	     data_out <= data_out_f;
	 when others =>
	     null;
    end case;

    ce(0)  <= cs and not( addr(14) ) and not( addr(13) ) and not( addr(12) ) and not( addr(11) );
    ce(1)  <= cs and not( addr(14) ) and not( addr(13) ) and not( addr(12) ) and      addr(11)  ;
    ce(2)  <= cs and not( addr(14) ) and not( addr(13) ) and      addr(12)   and not( addr(11) );
    ce(3)  <= cs and not( addr(14) ) and not( addr(13) ) and      addr(12)   and      addr(11)  ;
    ce(4)  <= cs and not( addr(14) ) and      addr(13)   and not( addr(12) ) and not( addr(11) );
    ce(5)  <= cs and not( addr(14) ) and      addr(13)   and not( addr(12) ) and      addr(11)  ;
    ce(6)  <= cs and not( addr(14) ) and      addr(13)   and      addr(12)   and not( addr(11) );
    ce(7)  <= cs and not( addr(14) ) and      addr(13)   and      addr(12)   and      addr(11)  ;
    ce(8)  <= cs and      addr(14)   and not( addr(13) ) and not( addr(12) ) and not( addr(11) );
    ce(9)  <= cs and      addr(14)   and not( addr(13) ) and not( addr(12) ) and      addr(11)  ;
    ce(10) <= cs and      addr(14)   and not( addr(13) ) and      addr(12)   and not( addr(11) );
    ce(11) <= cs and      addr(14)   and not( addr(13) ) and      addr(12)   and      addr(11)  ;
    ce(12) <= cs and      addr(14)   and      addr(13)   and not( addr(12) ) and not( addr(11) );
    ce(13) <= cs and      addr(14)   and      addr(13)   and not( addr(12) ) and      addr(11)  ;
    ce(14) <= cs and      addr(14)   and      addr(13)   and      addr(12)   and not( addr(11) );
    ce(15) <= cs and      addr(14)   and      addr(13)   and      addr(12)   and      addr(11)  ;

end process;

end architecture rtl;

