--===========================================================================--
--                                                                           --
--  sys09bug_s3e_rom2k_b16.vhd - Sys09bug monitor ROM for the Spartan 3E500  -- 
--                                                                           --
--===========================================================================--
--
--  File name      : sys09bug_s3e_rom2k_b16.vhd
--
--  Entity name    : mon_rom
--
--  Purpose        : Implements 2K Monitor ROM for System09
--                   using 1 x Spartan 3E RAMB16_S9 block ram
--                   Used in the Digilent Spartan 3E500 System09 design
--                  
--  Dependencies   : ieee.Std_Logic_1164
--                   ieee.std_logic_arith
--                   unisim.vcomponents
--
--  Uses           : RAMB16_S9
--
--  Author         : John E. Kent
--
--  Email          : dilbert57@opencores.org      
--
--  Web            : http://opencores.org/project,system09
--
--
--  Copyright (C) 2008 - 2010 John Kent
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--===========================================================================--
--                                                                           --
--                              Revision  History                            --
--                                                                           --
--===========================================================================--
--
-- Version Author      Date          Changes
-- 0.1     John Kent   2008-01-08    Initial Version
-- 0.2     John Kent   2010-09-14    Added Header
--                                   renamed rdata & wdata to data_out & data_in
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.vcomponents.all;

entity mon_rom is
    Port (
       clk      : in  std_logic;
       rst      : in  std_logic;
       cs       : in  std_logic;
       addr     : in  std_logic_vector (10 downto 0);
       rw       : in  std_logic;
       data_in  : in  std_logic_vector (7 downto 0);
       data_out : out std_logic_vector (7 downto 0)
    );
end mon_rom;

architecture rtl of mon_rom is

signal we : std_logic;
signal dp : std_logic;

begin

  MON_ROM : RAMB16_S9
    generic map ( 
         INIT_00 => x"A780A610C6C07F8E1060FE8EE0FE1FFB23FB94FBCFFCBAFC9CFCA2FC4BF814F8",
         INIT_01 => x"17431FE4A7D0866AAFDD8C30FB265AE26F0CC6450117D07FBF00E08EF9265AA0",
         INIT_02 => x"092C2081891FF1270D817F844E0417CE021794FE8EDE01174C031770FE8EA404",
         INIT_03 => x"FE8C02300F2780E12AFE8E20C0022F60C15E0417630417408B981F6A04175E86",
         INIT_04 => x"1F8002179CFE8E121F2D298603173B341FBC2094ADC0200B031796FE8EF52660",
         INIT_05 => x"17275E81DD271881E127088111287903171E0417C00317A4A6260417C0031721",
         INIT_06 => x"321FBD0217BE203F31C2202131FC03173F86FF03170827A4A1A4A7390F260D81",
         INIT_07 => x"F0C4201F0634F0C41000C3101F390124E1AC2034062926031705201F30C07F8E",
         INIT_08 => x"10C6AD0317490317E4AE0902179CFE8E10343962320327B103170527E4AC011F",
         INIT_09 => x"03172E8602237E810425208180A610C6E1AE9D0317F5265AA5031747031780A6",
         INIT_0a => x"273F8184A60F2710355B8DFFFF8E10341A24C07F8C1E29D20217BC20EE265A8E",
         INIT_0b => x"431F39FB265A1E8D08C6D37F8E105D03163F866003173984A73F86A4AFA0A709",
         INIT_0c => x"A60A24C07F8C21AEB3FE16ED7FBF00008E6302170C8D4AAF04272C8D1F304AAE",
         INIT_0d => x"265A0427A1ACA0A608C6D37F8E1039A0A7A0A7A0A7FF8684A7A4A604263F8184",
         INIT_0e => x"7FBFE7F98EEB7FBFC07FBEED7FBF14294B02170003171C29710117393D3139F7",
         INIT_0f => x"27ED7FBE24273F8184A64AAEFE011770E0B671E0B73686431F392020450017C0",
         INIT_10 => x"3B71E0B73F8673E0B7368670E0B671E0B7368670E0B70D86341FED7FBF1F301F",
         INIT_11 => x"B7368672E0B7008670E0B7FF8673E0B73A8671E0B7328622FE16C07FBFEB7FBE",
         INIT_12 => x"81380217D27F7F7602171186E8FCBD8435FD265A20C604343973E0B73E8671E0",
         INIT_13 => x"E0EBE0E610342129A3011726290234BA0117F12631813D273981310217F92653",
         INIT_14 => x"FFC102355FEB2080A70527E46AE0EB02340C290435A001170434E46AE46AE4EB",
         INIT_15 => x"02161386D27F73DE0117E101177801177B01177E01178101172802173F86BA27",
         INIT_16 => x"062762A3E4ECF501171286E8FCBDE4AF0130492562AC4D2930344A0117E26F0E",
         INIT_17 => x"63EB62EB68011762AE750117981F03CB2F0017DDFE8E64E720C6022320008310",
         INIT_18 => x"8D396532B301171486C326E4AC62AF5B0117981F53F526646A65011780A684EB",
         INIT_19 => x"AF0229F68DF28D910017E50016F800169D011690356900178EFE8E1034712002",
         INIT_1a => x"0229D58DD18D5E8D3946AF0229E08DDC8D728D3948AF0229EB8DE78D618D394A",
         INIT_1b => x"29B18DB08D588D3942A70229BC8DBB8D6C8D3943A70229C78DC68D498D3944AF",
         INIT_1c => x"F48DA0FE8E39F726048180A63B011739C4A7808A0429A68DA58D5F8D3941A702",
         INIT_1d => x"2044AED78DB8FE8EB4001643A6E18DBEFE8EF42048AEEA8DACFE8EBF0016311F",
         INIT_1e => x"8DC9FE8ED92041A6BC8DC4FE8ECF204AAEC58DA6FE8ED82046AECE8DB2FE8EE1",
         INIT_1f => x"B88DB08DA98DA18D27FF179CFE8E900016D5FE8EC4A6AA8DCEFE8ED02042A6B3",
         INIT_20 => x"1F42290E8DB400172D86121F4D29098DD520CE8DC78DC08D17FF179CFE8EBF8D",
         INIT_21 => x"578D39E0AB04342829078D891F484848483229118D903561A710343C29088D01",
         INIT_22 => x"578003226681072561813937800322468112254181393080032239811D253081",
         INIT_23 => x"078B022F3981308B0F840235048D4444444402340235028D0235103439021A39",
         INIT_24 => x"7F84048D0627D27F7D8235F1265A3B8D3F8D2D860225E46880A608C602344D20",
         INIT_25 => x"D07F9FA60234903501A6EE27018584A620E08E0926018584A6D07FBE10342D20",
         INIT_26 => x"F6260885FA27028584A6D07FBE1234498D2086008D8235018520E0B605260185",
         INIT_27 => x"00CC30E08E39D27FB7FF86016D84A7518684A70386D07FBE138D903501A70235",
         INIT_28 => x"7D30E08E16345986028D1B86F27F7F01E702C6F17FFD04E703E702A7EF7FFD00",
         INIT_29 => x"815A271B81342708819635AF001784A70520098D042420810D20608D0427F27F",
         INIT_2a => x"C15CEF7FFC45260A810F270B8124270C81890027100D81382716817C0027101A",
         INIT_2b => x"20212750814CEF7FB662204A2C27EF7FB66D205A34275DEF7FFC8F0016792619",
         INIT_2c => x"F27F7F39F27FB704263D81312754816E27598114273DC1F27FF656200000CC58",
         INIT_2d => x"20E12218C120C0F17F7FF17FF6ED224F812080F27F7F39F17FB70426F17F7D39",
         INIT_2e => x"A7EF7FFDF07FF64F39F27F7FF726508102A74C84E720C6EF7FB6168D0000CC1B",
         INIT_2f => x"F604E75F012519C15C04E6E78D5AEA2619C15C4FF02650814CEF7FFC3903E702",
         INIT_30 => x"E4205F03E7F07FF7082719C15CF07FF6F42650C15C84A702E7EF7FF72086EF7F",
         INIT_31 => x"1958FB1842FB1536FB1063FB0484FB036EFB0279FB0139F27FF702E7EF7FF75F",
         INIT_32 => x"C5F95472F958DBF853F2FB5292F84DC1FA5051FA4C8FF847E7F84546F9424DFB",
         INIT_33 => x"4F462047554239305359530000000A0DFFFFFFFF7EF991F891F891F891F87EF9",
         INIT_34 => x"04202D20043F54414857043E040000000A0D4B04202D2048544E5953444D2052",
         INIT_35 => x"2020043D58492020043D59492020043D53552020043D43502020043D50532020",
         INIT_36 => x"04315343565A4E4948464504203A43432020043D422020043D412020043D5044",
         INIT_37 => x"7F9F6EC87F9F6EC67F9F6EC47F9F6EC07F9F6E27F916D27FF7535FC07FCE1039",
         INIT_38 => x"AEC4EC10340822CE7FBC8B300F27FFFF8CCC7FBE49584F4AAF80E64AAE431FCA",
         INIT_39 => x"000000000000000000000000000000000000000000C27F9F6E42EE1F37F16E44",
         INIT_3a => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3b => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3c => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3d => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3e => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3f => x"E1FEEDFEFDFEF9FEF5FEF1FE01FFEDFE00000000000000000000000000000000"
    )

    port map (
	  do   => data_out,
	  dop(0) => dp,
	  addr => addr,
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp,
	  en   => cs,
	  ssr  => rst,
	  we   => we
	);

my_sbug : process ( rw )
begin
	 we    <= not rw;
end process;

end architecture rtl;

