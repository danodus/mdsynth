--===========================================================================--
--                                                                           --
--  sys09bug_s3e_rom2k_b16.vhd - Sys09bug monitor ROM for the Spartan 3E500  -- 
--                                                                           --
--===========================================================================--
--
--  File name      : sys09bug_s3e_rom2k_b16.vhd
--
--  Entity name    : mon_rom
--
--  Purpose        : Implements 2K Monitor ROM for System09
--                   using 1 x Spartan 3E RAMB16_S9 block ram
--                   Used in the Digilent Spartan 3E500 System09 design
--                  
--  Dependencies   : ieee.Std_Logic_1164
--                   ieee.std_logic_arith
--                   unisim.vcomponents
--
--  Uses           : RAMB16_S9
--
--  Author         : John E. Kent
--
--  Email          : dilbert57@opencores.org      
--
--  Web            : http://opencores.org/project,system09
--
--
--  Copyright (C) 2008 - 2010 John Kent
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--===========================================================================--
--                                                                           --
--                              Revision  History                            --
--                                                                           --
--===========================================================================--
--
-- Version Author      Date          Changes
-- 0.1     John Kent   2008-01-08    Initial Version
-- 0.2     John Kent   2010-09-14    Added Header
--                                   renamed rdata & wdata to data_out & data_in
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
	use unisim.vcomponents.all;

entity mon_rom is
    Port (
       clk      : in  std_logic;
       rst      : in  std_logic;
       cs       : in  std_logic;
       addr     : in  std_logic_vector (10 downto 0);
       rw       : in  std_logic;
       data_in  : in  std_logic_vector (7 downto 0);
       data_out : out std_logic_vector (7 downto 0)
    );
end mon_rom;

architecture rtl of mon_rom is

signal we : std_logic;
signal dp : std_logic;

begin

  MON_ROM : RAMB16_S9
    generic map ( 
         INIT_00 => x"A780A610C6C07F8E104EFE8ECEFE0DFB11FB82FBBDFCA8FC8AFC90FC4BF814F8",
         INIT_01 => x"17431FE4A7D0866AAFDD8C30FB265AE26F0CC6450117D07FBF00E08EF9265AA0",
         INIT_02 => x"092C2081891FF1270D817F843C0417BC021782FE8EDE01173A03175EFE8E9204",
         INIT_03 => x"FE8C02300F2780E118FE8E20C0022F60C14C0417510417408B981F5804175E86",
         INIT_04 => x"1F6E02178AFE8E121F2D297403173B341FBC2094ADC020F9021784FE8EF5264E",
         INIT_05 => x"17275E81DD271881E127088111286703170C0417AE0317A4A6140417AE031721",
         INIT_06 => x"321FAB0217BE203F31C2202131EA03173F86ED03170827A4A1A4A7390F260D81",
         INIT_07 => x"F0C4201F0634F0C41000C3101F390124E1AC2034062914031705201F30C07F8E",
         INIT_08 => x"10C69B0317370317E4AEF701178AFE8E103439623203279F03170527E4AC011F",
         INIT_09 => x"03172E8602237E810425208180A610C6E1AE8B0317F5265A93031735031780A6",
         INIT_0a => x"273F8184A60F2710355B8DFFFF8E10341A24C07F8C1E29C00217BC20EE265A7C",
         INIT_0b => x"431F39FB265A1E8D08C6D37F8E104B03163F864E03173984A73F86A4AFA0A709",
         INIT_0c => x"A60A24C07F8C21AEB3FE16ED7FBF00008E5102170C8D4AAF04272C8D1F304AAE",
         INIT_0d => x"265A0427A1ACA0A608C6D37F8E1039A0A7A0A7A0A7FF8684A7A4A604263F8184",
         INIT_0e => x"7FBFE7F98EEB7FBFC07FBEED7FBF1429390217EE02171C295F0117393D3139F7",
         INIT_0f => x"27ED7FBE24273F8184A64AAEEC011770E0B671E0B73686431F392020450017C0",
         INIT_10 => x"3B71E0B73F8673E0B7368670E0B671E0B7368670E0B70D86341FED7FBF1F301F",
         INIT_11 => x"B7368672E0B7008670E0B7FF8673E0B73A8671E0B7328622FE16C07FBFEB7FBE",
         INIT_12 => x"81260217D27F7F6402171186D6FCBD8435FD265A20C604343973E0B73E8671E0",
         INIT_13 => x"E0EBE0E61034212991011726290234A80117F12631813D2739811F0217F92653",
         INIT_14 => x"FFC102355FEB2080A70527E46AE0EB02340C2904358E01170434E46AE46AE4EB",
         INIT_15 => x"E4AF0130492562AC4D2930344A0117E26F0E02161386D27F731602173F86BA27",
         INIT_16 => x"03CB2F0017CBFE8E64E720C6022320008310062762A3E4ECF501171286D6FCBD",
         INIT_17 => x"AF5B0117981F53F526646A65011780A684EB63EB62EB68011762AE750117981F",
         INIT_18 => x"00169D011690356900177CFE8E10347120028D396532B301171486C326E4AC62",
         INIT_19 => x"8DDC8D728D3948AF0229EB8DE78D618D394AAF0229F68DF28D910017E50016F8",
         INIT_1a => x"BB8D6C8D3943A70229C78DC68D498D3944AF0229D58DD18D5E8D3946AF0229E0",
         INIT_1b => x"1739C4A7808A0429A68DA58D5F8D3941A70229B18DB08D588D3942A70229BC8D",
         INIT_1c => x"8DACFE8EF42048AEEA8D9AFE8EBF0016311FF48D8EFE8E39F726048180A63B01",
         INIT_1d => x"204AAEC58D94FE8ED82046AECE8DA0FE8EE12044AED78DA6FE8EB4001643A6E1",
         INIT_1e => x"900016C3FE8EC4A6AA8DBCFE8ED02042A6B38DB7FE8ED92041A6BC8DB2FE8ECF",
         INIT_1f => x"098DD520CE8DC78DC08D17FF178AFE8EBF8DB88DB08DA98DA18D27FF178AFE8E",
         INIT_20 => x"4848483229118D903561A710343C29088D011F42290E8DB400172D86121F4D29",
         INIT_21 => x"22468112254181393080032239811D253081578D39E0AB04342829078D891F48",
         INIT_22 => x"4444444402340235028D0235103439021A395780032266810725618139378003",
         INIT_23 => x"3B8D3F8D2D860225E46880A608C602344D20078B022F3981308B0F840235048D",
         INIT_24 => x"84A620E08E0926018584A6D07FBE10342D207F84048D0627D27F7D8235F1265A",
         INIT_25 => x"34498D2086008D8235018520E0B605260185D07F9FA60234903501A6EE270185",
         INIT_26 => x"A7518684A70386D07FBE138D903501A70235F6260885FA27028584A6D07FBE12",
         INIT_27 => x"7F01E702C6F17FFD04E703E702A7EF7FFD0000CC30E08E39D27FB7FF86016D84",
         INIT_28 => x"84A70520098D042420810D20608D0427F27F7D30E08E16345986028D1B86F27F",
         INIT_29 => x"270C81890027100D81382716817C0027101A815A271B81342708819635AF0017",
         INIT_2a => x"EF7FB66D205A34275DEF7FFC8F0016792619C15CEF7FFC45260A810F270B8124",
         INIT_2b => x"816E27598114273DC1F27FF656200000CC5820212750814CEF7FB662204A2C27",
         INIT_2c => x"224F812080F27F7F39F17FB70426F17F7D39F27F7F39F27FB704263D81312754",
         INIT_2d => x"508102A74C84E720C6EF7FB6168D0000CC1B20E12218C120C0F17F7FF17FF6ED",
         INIT_2e => x"EA2619C15C4FF02650814CEF7FFC3903E702A7EF7FFDF07FF64F39F27F7FF726",
         INIT_2f => x"7FF6F42650C15C84A702E7EF7FF72086EF7FF604E75F012519C15C04E6E78D5A",
         INIT_30 => x"FB035CFB0267FB0139F27FF702E7EF7FF75FE4205F03E7F07FF7082719C15CF0",
         INIT_31 => x"4DAFFA5051FA4C8FF847E7F84546F9423BFB1946FB1830FB1524FB1051FB0472",
         INIT_32 => x"0A0DFFFFFFFF7EF991F891F891F891F87EF9C5F95472F958DBF853E0FB5292F8",
         INIT_33 => x"00000A0D4B04202D2048544E5953444D20524F46204755423930535953000000",
         INIT_34 => x"043D53552020043D43502020043D5053202004202D20043F54414857043E0400",
         INIT_35 => x"43432020043D422020043D412020043D50442020043D58492020043D59492020",
         INIT_36 => x"6EC07F9F6E39F916D27FF7535FC07FCE103904315343565A4E4948464504203A",
         INIT_37 => x"FFFF8CCC7FBE49584F4AAF80E64AAE431FCA7F9F6EC87F9F6EC67F9F6EC47F9F",
         INIT_38 => x"00000000000000C27F9F6E42EE1F37F16E44AEC4EC10340822CE7FBC8B300F27",
         INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3a => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3b => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3c => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3d => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3e => x"0000000000000000000000000000000000000000000000000000000000000000",
         INIT_3f => x"CFFEDBFEEBFEE7FEE3FEDFFEEFFEDBFE00000000000000000000000000000000"
    )

    port map (
	  do   => data_out,
	  dop(0) => dp,
	  addr => addr,
	  clk  => clk,
     di   => data_in,
	  dip(0) => dp,
	  en   => cs,
	  ssr  => rst,
	  we   => we
	);

my_sbug : process ( rw )
begin
	 we    <= not rw;
end process;

end architecture rtl;

